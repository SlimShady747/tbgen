// Generatated test bench (sample tbgen.py template)
`default_nettype none
%%%TIMESCALE%%%
%%%HEAD%%%
%%%WIRES%%%
%%%UUT%%% (
%%%ARGS%%% );
%%%PERIOD%%%
%%%CLOCK%%%
initial begin
%%%DUMP%%%
end
initial begin
%%%RESET%%%
end
// Include your custom changes in the included file
%%%INCLUDE%%%

endmodule
